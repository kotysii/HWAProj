`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 01.12.2019 18:44:41
// Design Name: 
// Module Name: APractice
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module APractice(input[3:0] in, output[3:0] out);
    out[2] != in[2]
    out[1] != in[1]
    out[0] != in[0]
    
endmodule
