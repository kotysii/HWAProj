`timescale 1ns / 1ps

module APractice(input[3:0] in, output[3:0] out);

assign 
    
endmodule
